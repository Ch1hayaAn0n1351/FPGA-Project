`timescale 1ns/1ps
module vga_pic(
    input wire vga_clk ,
    input wire sys_rst_n ,
    input wire [9:0] pix_x ,
    input wire [9:0] pix_y ,
    output reg [15:0] pix_data
);

parameter H_VALID   = 10'd640;
parameter V_VALID   = 10'd480;
parameter CHAR_W    = 10'd32;
parameter CHAR_H    = 10'd32;
parameter BYTE_PER_ROW = 4;
parameter RED       = 16'hF800;
parameter BLACK     = 16'h0000;

localparam TOTAL_CHAR_W = 4 * CHAR_W;
localparam START_X = (H_VALID - TOTAL_CHAR_W) / 2;
localparam START_Y = (V_VALID - CHAR_H) / 2;

reg [7:0] m_bitmap [31:0][BYTE_PER_ROW-1:0];
reg [7:0] u_bitmap [31:0][BYTE_PER_ROW-1:0];
reg [7:0] s_bitmap [31:0][BYTE_PER_ROW-1:0];
reg [7:0] t_bitmap [31:0][BYTE_PER_ROW-1:0];

initial begin
    for (integer i = 0; i < 32; i = i + 1) begin
        m_bitmap[i][0] = {0x00,0x00,0x00,0x00,0x00,0x00,0xf8,0x78,0x78,0x78,0x7c,0x7c,0x7c,0x7c,0x7e,0x7e,0x7e,0x6e,0x6e,0x6f,0x6f,0x6f,0x67,0x67,0x67,0x67,0x73,0xfb,0x00,0x00,0x00,0x00}[i];
        m_bitmap[i][1] = {0x00,0x00,0x00,0x00,0x00,0x00,0x1f,0x3e,0x3e,0x3e,0x3e,0x7e,0x7e,0x7e,0x7e,0x7e,0xfe,0xfe,0xfe,0xde,0xde,0xde,0xde,0x9e,0x9e,0x9e,0x9e,0x7f,0x00,0x00,0x00,0x00}[i];
        m_bitmap[i][2] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
        m_bitmap[i][3] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
    end

    for (integer i = 0; i < 32; i = i + 1) begin
        u_bitmap[i][0] = {0x00,0x00,0x00,0x00,0x00,0x00,0xfe,0x7c,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x78,0x38,0x38,0x3c,0x1f,0x0f,0x00,0x00,0x00,0x00}[i];
        u_bitmap[i][1] = {0x00,0x00,0x00,0x00,0x00,0x00,0x3f,0x1e,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x0c,0x1c,0x3c,0xf8,0xf0,0x00,0x00,0x00,0x00}[i];
        u_bitmap[i][2] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
        u_bitmap[i][3] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
    end

    for (integer i = 0; i < 32; i = i + 1) begin
        s_bitmap[i][0] = {0x00,0x00,0x00,0x00,0x00,0x00,0x1f,0x3e,0x38,0x70,0x70,0x70,0x78,0x7c,0x3f,0x3f,0x0f,0x03,0x00,0x00,0x00,0x60,0x60,0x70,0x70,0x78,0x7f,0x7f,0x00,0x00,0x00,0x00}[i];
        s_bitmap[i][1] = {0x00,0x00,0x00,0x00,0x00,0x00,0xfc,0xfc,0x3c,0x1c,0x1c,0x0c,0x00,0x00,0x00,0xc0,0xf0,0xf8,0xfc,0x3c,0x1e,0x1e,0x0e,0x1e,0x1e,0x3c,0xf8,0xf0,0x00,0x00,0x00,0x00}[i];
        s_bitmap[i][2] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
        s_bitmap[i][3] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
    end

    for (integer i = 0; i < 32; i = i + 1) begin
        t_bitmap[i][0] = {0x00,0x00,0x00,0x00,0x00,0x00,0x7f,0x7b,0x73,0xe3,0xe3,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x03,0x0f,0x00,0x00,0x00,0x00}[i];
        t_bitmap[i][1] = {0x00,0x00,0x00,0x00,0x00,0x00,0xfe,0xde,0xce,0xc6,0xc7,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xc0,0xf0,0x00,0x00,0x00,0x00}[i];
        t_bitmap[i][2] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
        t_bitmap[i][3] = {0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00}[i];
    end
end

always @(posedge vga_clk or negedge sys_rst_n) begin
    if (!sys_rst_n) begin
        pix_data <= BLACK;
    end else begin
        if ((pix_y >= START_Y) && (pix_y < START_Y + CHAR_H) && 
            (pix_x >= START_X) && (pix_x < START_X + TOTAL_CHAR_W)) begin
            
            reg [4:0] char_y;
            reg [6:0] char_x;
            reg [1:0] byte_idx;
            reg [2:0] bit_idx;
            
            char_y = pix_y - START_Y;
            char_x = pix_x - START_X;

            if (char_x < CHAR_W) begin
                byte_idx = char_x[4:3];
                bit_idx  = char_x[2:0];
                pix_data = (m_bitmap[char_y][byte_idx][7 - bit_idx]) ? RED : BLACK;
            end else if (char_x < 2*CHAR_W) begin
                char_x = char_x - CHAR_W;
                byte_idx = char_x[4:3];
                bit_idx  = char_x[2:0];
                pix_data = (u_bitmap[char_y][byte_idx][7 - bit_idx]) ? RED : BLACK;
            end else if (char_x < 3*CHAR_W) begin
                char_x = char_x - 2*CHAR_W;
                byte_idx = char_x[4:3];
                bit_idx  = char_x[2:0];
                pix_data = (s_bitmap[char_y][byte_idx][7 - bit_idx]) ? RED : BLACK;
            end else begin
                char_x = char_x - 3*CHAR_W;
                byte_idx = char_x[4:3];
                bit_idx  = char_x[2:0];
                pix_data = (t_bitmap[char_y][byte_idx][7 - bit_idx]) ? RED : BLACK;
            end
        end else begin
            pix_data <= BLACK;
        end
    end
end

endmodule
endmodule
